// Listing 14.3
/******************************************************************
* Mark1 Mod:
* - invert reset signal
********************************************************************/
module font_test_top
   (
    input wire clk, reset,
    output wire hsync, vsync,
    output wire [2:0] rgb
   );

   // signal declaration
   wire [9:0] pixel_x, pixel_y;
   wire video_on, pixel_tick;
   reg [2:0] rgb_reg;
   wire [2:0] rgb_next;
	wire nreset;	//invert reset signal
	
	assign nreset = ~reset;

   // body
   // instantiate vga sync circuit
   vga_sync vsync_unit
      (	.clk(clk), 
			.reset(nreset), 
			.hsync(hsync), 
			.vsync(vsync),
			.video_on(video_on), 
			.p_tick(pixel_tick),
			.pixel_x(pixel_x), 
			.pixel_y(pixel_y)
		);
   // font generation circuit
   font_test_gen font_gen_unit
      (	.clk(clk), 
			.video_on(video_on), 
			.pixel_x(pixel_x),
			.pixel_y(pixel_y), 
			.rgb_text(rgb_next)
		);
   // rgb buffer
   always @(posedge clk)
      if (pixel_tick)
         rgb_reg <= rgb_next;
   // output
   assign rgb = rgb_reg;

endmodule

