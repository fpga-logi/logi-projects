----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    14:14:22 06/21/2012 
-- Design Name: 
-- Module Name:    spartcam_beaglebone - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

library work ;
use work.utils_pack.all ;
use work.peripheral_pack.all ;
use work.interface_pack.all ;
use work.conf_pack.all ;
use work.filter_pack.all ;
use work.image_pack.all ;
use work.blob_pack.all ;
use work.classifier_pack.all ;
use work.primitive_pack.all ;
-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
library UNISIM;
use UNISIM.VComponents.all;

entity mark1_rpi_blob_tracking is
port( OSC_FPGA : in std_logic;

		--onboard
		PB, DIP_SW : in std_logic_vector(3 downto 0);
		LED : out std_logic_vector(7 downto 0);	
		
			--PMOD
		PMOD4_6, PMOD4_2  : inout std_logic ; -- used as SCL, SDA
		PMOD4_0, PMOD4_3 : out std_logic ; -- used as reset and xclk 
		PMOD4_7, PMOD4_1, PMOD4_5, PMOD4_4 : in std_logic ; -- used as pclk, href, vsync
		PMOD3 : in std_logic_vector(7 downto 0); -- used as cam data
		
		
		--i2c
		SYS_I2C_SCL, SYS_I2C_SDA : inout std_logic ;
		
		--spi
		SYS_SPI_SCK, SYS_SPI_SS, SYS_SPI_MOSI : in std_logic ;
		SYS_SPI_MISO : out std_logic 
);
end mark1_rpi_blob_tracking;

architecture Behavioral of mark1_rpi_blob_tracking is

	COMPONENT clock_gen
	PORT(
		CLK_IN1 : IN std_logic;          
		CLK_OUT1 : OUT std_logic;
		CLK_OUT2 : OUT std_logic;
		CLK_OUT3 : OUT std_logic;
		LOCKED : OUT std_logic
		);
	END COMPONENT;

	
	signal clk_sys, clk_100, clk_24, clk_locked : std_logic ;
	signal resetn , sys_resetn : std_logic ;
	
	signal counter_output : std_logic_vector(31 downto 0);
	signal fifo_output : std_logic_vector(15 downto 0);
	signal fifo_input : std_logic_vector(15 downto 0);
	signal color_lut_data_out : std_logic_vector(15 downto 0);
	signal image_fifo_wr : std_logic ;
	signal blob_fifo_input : std_logic_vector(15 downto 0);
	signal bus_blob_fifo_out : std_logic_vector(15 downto 0);
	signal blob_fifo_wr, cs_blob_fifo : std_logic ;
	signal bus_data_in, bus_data_out : std_logic_vector(15 downto 0);
	signal bus_fifo_out, bus_latch_out : std_logic_vector(15 downto 0);
	signal bus_addr : std_logic_vector(15 downto 0);
	signal bus_wr, bus_rd, bus_cs : std_logic ;
	signal cs_image_fifo, cs_color_lut : std_logic ;
	signal color_index : std_logic_vector(15 downto 0);
	
	signal cam_data : std_logic_vector(7 downto 0);
	signal cam_sioc, cam_siod : std_logic ;
	signal cam_xclk, cam_pclk, cam_vsync, cam_href, cam_reset : std_logic ;
	
	signal rom_addr : std_logic_vector(7 downto 0);
	signal rom_data : std_logic_vector(15 downto 0);
	
	signal pixel_y_from_interface, pixel_u_from_interface, pixel_v_from_interface : std_logic_vector(7 downto 0);
	signal pxclk_from_interface, href_from_interface, vsync_from_interface : std_logic ;
	signal pixel_from_bin : std_logic_vector(7 downto 0);
	signal pxclk_from_bin, href_from_bin, vsync_from_bin : std_logic ;
	signal pixel_from_erode : std_logic_vector(7 downto 0);
	signal pxclk_from_erode, href_from_erode, vsync_from_erode : std_logic ;
	signal pixel_low_thresh, pixel_high_thresh : std_logic_vector(7 downto 0);
	
	
	signal output_pxclk, output_href , output_vsync : std_logic ;
	signal output_pixel : std_logic_vector(7 downto 0);
	signal hsync_rising_edge, vsync_rising_edge, pxclk_rising_edge, hsync_old, vsync_old, pxclk_old, write_pixel_old : std_logic ;
	signal pixel_buffer : std_logic_vector(15 downto 0);	
	signal pixel_count :std_logic_vector(7 downto 0);
	signal write_pixel : std_logic ;
	
	signal color_lut_out : std_logic_vector(7 downto 0);
	
	for all : yuv_register_rom use entity work.yuv_register_rom(ov7725_qvga);
begin
	
	resetn <= PB(0) ;
	sys_clocks_gen: clock_gen 
	PORT MAP(
		CLK_IN1 => OSC_FPGA,
		CLK_OUT1 => clk_100,
		CLK_OUT2 => clk_24,
		CLK_OUT3 => clk_sys, --120Mhz system clock
		LOCKED => clk_locked
	);


	reset0: reset_generator 
	generic map(HOLD_0 => 1000)
	port map(clk => clk_sys, 
		resetn => resetn ,
		resetn_0 => sys_resetn
	 );


divider : simple_counter 
	 generic map(NBIT => 32)
    port map( clk => clk_sys, 
           resetn => sys_resetn, 
           sraz => '0',
           en => '1',
			  load => '0' ,
			  E => X"00000000",
			  Q => counter_output
			  );
LED(0) <= counter_output(24);
LED(1) <= cam_vsync;
LED(2) <= cam_href;
LED(3) <= not cs_blob_fifo ;
LED(4) <= not cs_image_fifo;
LED(7 downto 5) <= counter_output(27 downto 25);


mem_interface0 : spi2ad_bus
generic map(ADDR_WIDTH => 16 , DATA_WIDTH =>  16)
port map(clk => clk_sys ,
	  resetn => sys_resetn ,
	  mosi => SYS_SPI_MOSI,
	  miso => SYS_SPI_MISO,
	  sck => SYS_SPI_SCK,
	  ss => SYS_SPI_SS,
	  data_bus_out	=> bus_data_out,
	  data_bus_in	=> bus_data_in ,
	  addr_bus	=> bus_addr, 
	  wr => bus_wr , rd => bus_rd 
);

cs_image_fifo <= '1' when bus_addr(15 downto 3) = "0000000000000" else
			  '0' ;

cs_blob_fifo <= '1' when bus_addr(15 downto 3) = "0000000000001" else
			  '0' ;
			  
cs_color_lut <= '1' when bus_addr(15 downto 12) = "0001" else
			  '0' ;

bus_data_in <= bus_fifo_out when cs_image_fifo = '1' else
					bus_blob_fifo_out when cs_blob_fifo = '1' else
					color_lut_data_out when cs_color_lut = '1' else
					(others => '1');

bi_fifo0 : fifo_peripheral 
		generic map(ADDR_WIDTH => 16,WIDTH => 16, SIZE => 4096, BURST_SIZE => 4)
		port map(
			clk => clk_sys,
			resetn => sys_resetn,
			addr_bus => bus_addr,
			wr_bus => bus_wr,
			rd_bus => bus_rd,
			cs_bus => cs_image_fifo,
			wrB => image_fifo_wr,
			rdA => '0',
			data_bus_in => bus_data_out,
			data_bus_out => bus_fifo_out,
			inputB => fifo_input, 
			outputA => open,
			emptyA => open,
			fullA => open,
			emptyB => open,
			fullB => open,
			burst_available_B => open
		);

fifo_blobs : fifo_peripheral 
		generic map(ADDR_WIDTH => 16,
						WIDTH => 16, 
						SIZE => 1024, 
						BURST_SIZE => 4,
						SYNC_LOGIC_INTERFACE => true)
		port map(
			clk => clk_sys,
			resetn => sys_resetn,
			addr_bus => bus_addr,
			wr_bus => bus_wr,
			rd_bus => bus_rd,
			cs_bus => cs_blob_fifo,
			wrB => blob_fifo_wr,
			rdA => '0',
			data_bus_in => bus_data_out,
			data_bus_out => bus_blob_fifo_out,
			inputB => blob_fifo_input, 
			outputA => open,
			emptyA => open,
			fullA => open,
			emptyB => open,
			fullB => open,
			burst_available_B => open
		);		
 
 conf_rom : yuv_register_rom
	port map(
	   clk => clk_sys, en => '1' ,
 		data => rom_data,
 		addr => rom_addr
	); 
 
 camera_conf_block : i2c_conf 
	generic map(ADD_WIDTH => 8 , SLAVE_ADD => "0100001")
	port map(
		clock => clk_sys, 
		resetn => sys_resetn ,		
 		i2c_clk => clk_24 ,
		scl => PMOD4_6,
 		sda => PMOD4_2, 
		reg_addr => rom_addr ,
		reg_data => rom_data
	);	
		
 camera0: yuv_camera_interface
		port map(clock => clk_sys,
					resetn => sys_resetn,
					pixel_data => cam_data, 
					pxclk => cam_pclk, href => cam_href, vsync => cam_vsync,
					pixel_clock_out => pxclk_from_interface, hsync_out => href_from_interface, vsync_out => vsync_from_interface,
					y_data => pixel_y_from_interface,
					u_data => pixel_u_from_interface,
					v_data => pixel_v_from_interface
					
		);	
		
	cam_xclk <= clk_24;
	PMOD4_3 <= cam_xclk ;
	--cam_data <= PMOD2 ;
	cam_data <= PMOD3(3) & PMOD3(7) & PMOD3(2) & PMOD3(6) & PMOD3(1) & PMOD3(5) & PMOD3(0) & PMOD3(4) ;
	cam_pclk <= PMOD4_7 ;
	cam_href <= PMOD4_1 ;
	cam_vsync <= PMOD4_5 ;
	PMOD4_0 <= cam_reset ;
	cam_reset <= resetn ;

classifier_lut : dpram_NxN	
	generic map(SIZE => 4096, NBIT => 2, ADDR_WIDTH => 12)
	port map(
 		clk => clk_sys ,
 		we =>  (bus_wr AND cs_color_lut),
 		
 		di => bus_data_out(1 downto 0), 
		a	=> bus_addr(11 downto 0),
 		dpra => color_index(11 downto 0),
		spo => color_lut_data_out(1 downto 0),
		dpo => color_lut_out(1 downto 0) 		
	); 

classification0 : color_classifier
port map( 		clk => clk_sys, 
 		resetn => sys_resetn ,
 		pixel_clock => pxclk_from_interface, hsync => href_from_interface, vsync => vsync_from_interface,
 		pixel_clock_out => pxclk_from_bin, hsync_out => href_from_bin, vsync_out => vsync_from_bin,
		pixel_y => pixel_y_from_interface,
		pixel_u => pixel_u_from_interface,
		pixel_v => pixel_v_from_interface,
		pixel_class => pixel_from_bin,
		
		color_index => color_index(11 downto 0),
		lut_in => color_lut_out
);


smooth0 : classifier_smoother 
generic map(WIDTH => 320, HEIGHT => 240)
port map(
 		clk => clk_sys, 
 		resetn => sys_resetn ,
 		pixel_clock => pxclk_from_bin, hsync => href_from_bin, vsync => vsync_from_bin,
 		pixel_clock_out => pxclk_from_erode, hsync_out => href_from_erode, vsync_out => vsync_from_erode,
 		pixel_data_in => pixel_from_bin,
 		pixel_data_out => pixel_from_erode
);


blob_tracker : blob_detection 
generic map(LINE_SIZE => 320)
port map(
 		clk => clk_sys, 
 		resetn => sys_resetn ,
 		pixel_clock => pxclk_from_erode, hsync => href_from_erode, vsync => vsync_from_erode,
		pixel_data_in => pixel_from_erode,
		blob_data => open,
		
		--memory_interface to copy results on vsync
		mem_addr => open,
		mem_data =>blob_fifo_input,
		mem_wr => blob_fifo_wr
);





output_pxclk <= pxclk_from_erode ;
output_href <= href_from_erode ;
output_vsync <= vsync_from_erode ;
output_pixel <= pixel_from_erode ;




--output_pxclk <= pxclk_from_interface ;
--output_href <= href_from_interface ;
--output_vsync <= vsync_from_interface ;
--output_pixel <= pixel_y_from_interface ;
	
--pix2fifo : pixel2fifo 
--port map(
--	clk => clk_sys, resetn => sys_resetn,
--	pixel_clock => output_pxclk, hsync => output_href, vsync => output_vsync,
--	pixel_data_in => output_pixel,
--	fifo_data => fifo_input, 
--	fifo_wr => image_fifo_wr 
--
--);


	
	process(clk_sys, sys_resetn)
begin
	if sys_resetn = '0' then
		vsync_old <= '0' ;
	elsif clk_sys'event and clk_sys = '1' then
		vsync_old <= output_vsync ;
	end if ;
end process ;
vsync_rising_edge <= (NOT vsync_old) and output_vsync ;

process(clk_sys, sys_resetn)
begin
	if sys_resetn = '0' then
		hsync_old <= '0' ;
	elsif clk_sys'event and clk_sys = '1' then
		hsync_old <= output_href ;
	end if ;
end process ;
hsync_rising_edge <= (NOT hsync_old) and output_href ;

process(clk_sys, sys_resetn)
begin
	if sys_resetn = '0' then
		pxclk_old <= '0' ;
	elsif clk_sys'event and clk_sys = '1' then
		pxclk_old <= output_pxclk ;
	end if ;
end process ;
pxclk_rising_edge <= (NOT pxclk_old) and output_pxclk ;

process(clk_sys, sys_resetn)
begin
	if sys_resetn = '0' then
		pixel_buffer(15 downto 0) <= (others => '0') ;
	elsif clk_sys'event and clk_sys = '1' then
		if hsync_rising_edge = '1' then
			pixel_buffer(15 downto 0) <= (others => '0') ;
		elsif pxclk_rising_edge = '1' then
			pixel_buffer(7 downto 0) <= pixel_buffer(15 downto 8) ;
			pixel_buffer(15 downto 8)  <= output_pixel ;
		end if ;
	end if ;
end process ;

process(clk_sys, sys_resetn)
begin
	if sys_resetn = '0' then
		pixel_count <= (others => '0'); 
	elsif clk_sys'event and clk_sys = '1' then
		if hsync_rising_edge = '1' then
			pixel_count <= (others => '0'); 
		elsif pxclk_rising_edge = '1'  and href_from_interface = '0' then
			pixel_count <= pixel_count + 1 ;
		end if ;
	end if ;
end process ;
write_pixel <= pixel_count(0);

process(clk_sys, sys_resetn)
begin
	if sys_resetn = '0' then
		write_pixel_old <= '0'; 
	elsif clk_sys'event and clk_sys = '1' then
		write_pixel_old <= write_pixel ;
	end if ;
end process ;


image_fifo_wr <= (write_pixel and (NOT write_pixel_old)) when output_vsync = '0' and output_href = '0' else
			   vsync_rising_edge when output_vsync = '1' else
				'0' ;
				
fifo_input <= (X"AA55") when vsync_rising_edge = '1' else
				  (pixel_buffer(15 downto 1) & '0') when pixel_buffer = X"AA55" else
				  pixel_buffer;

end Behavioral;

